.title KiCad schematic
.include "/usr/share/kicad/library/pspice.lib"
MU1 0 Net-_C1-Pad2_ Net-_C1-Pad1_ Net-_U1-Pad4_ Net-_U1-Pad5_ OPAMP
V1 Net-_U1-Pad4_ 0 dc 2.5
R2 Net-_C1-Pad1_ 0 100k
R1 Net-_C1-Pad1_ Net-_C1-Pad2_ 20
V2 0 Net-_U1-Pad5_ dc 2.5
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 1000p
I1 Net-_C1-Pad2_ 0 dc 20m
.end
